module main_decoder (
   op,
   branch,
   resultsrc,
   memwrite,
   alusrc,
   immsrc,
   regwrite,
   aluop
);



endmodule 